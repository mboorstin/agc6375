import GetPut::*;
import InterStage::*;
import Exec::*;

(* synthesize *)
module mkExecTest ();
    //


    //module to test
    //Exec exec <- mkExec();

    //test inputs
    Decode2Exec d2e;
    
endmodule

